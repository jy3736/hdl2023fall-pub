// write your module here