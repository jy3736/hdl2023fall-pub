module decode(
  input [3:0] din, 
  output reg odd, 
  output reg even,
  output reg zero
);

  // TODO: write your code here

endmodule