module router(
    input [7:0] a,
    input [7:0] b,
    input [1:0] sel,
    output [7:0] x,
    output [7:0] y
);

    // write your code here

endmodule
