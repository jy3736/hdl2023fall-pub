// write your module here
